// Author: Ujjval Raghavendra L

module top_module( input in, output out );
assign out = ~in;
endmodule
