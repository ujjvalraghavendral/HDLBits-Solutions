// Author: Ujjval Raghavendra L

module top_module(output zero);

endmodule
