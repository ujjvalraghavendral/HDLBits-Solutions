// Author: Ujjval Raghavendra L


module top_module (
    input c,
    input d,
    output [3:0] mux_in
); 
	// Split the truth table into four columns,
	assign mux_in[0] = c ? 1 : d;          // 1 mux:   c|d
	assign mux_in[1] = 0;                  // No muxes:  0
	assign mux_in[2] = d ? 0 : 1;          // 1 mux:    ~d
	assign mux_in[3] = c ? d : 0;          // 1 mux:   c&d

endmodule

